
module nios_system (
	clk_50_in_clk,
	reset_reset_n,
	clk_50_2_in_clk,
	reset_0_reset_n,
	clk_50_3_in_clk,
	reset_1_reset_n);	

	input		clk_50_in_clk;
	input		reset_reset_n;
	input		clk_50_2_in_clk;
	input		reset_0_reset_n;
	input		clk_50_3_in_clk;
	input		reset_1_reset_n;
endmodule


module avalon_timer_32b_qsys (
	clk_clk,
	reset_reset_n,
	avalon_timer_32b_external_interface_conduit0);	

	input		clk_clk;
	input		reset_reset_n;
	output		avalon_timer_32b_external_interface_conduit0;
endmodule

module top();
      avalon_timer_32b_qsys_tb tb ();
      test_program pgm ();
endmodule

// tangente_PWL_vhd.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module tangente_PWL_vhd (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

endmodule


module avalon_timer_32b_qsys (
	avalon_timer_32b_external_interface_conduit0,
	clk_clk,
	reset_reset_n);	

	output		avalon_timer_32b_external_interface_conduit0;
	input		clk_clk;
	input		reset_reset_n;
endmodule

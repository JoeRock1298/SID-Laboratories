
module nios_system (
	clock_50_clk,
	reset_reset_n,
	led_green_external_export);	

	input		clock_50_clk;
	input		reset_reset_n;
	output	[7:0]	led_green_external_export;
endmodule

// avalon_displays7seg_qsys_tb.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module avalon_displays7seg_qsys_tb (
	);

	wire        avalon_displays7seg_qsys_inst_clk_bfm_clk_clk;                          // avalon_displays7seg_qsys_inst_clk_bfm:clk -> [avalon_displays7seg_qsys_inst:clk_clk, avalon_displays7seg_qsys_inst_displays7seg_external_interface_bfm:clk, avalon_displays7seg_qsys_inst_reset_bfm:clk]
	wire  [6:0] avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit3; // avalon_displays7seg_qsys_inst:displays7seg_external_interface_conduit3 -> avalon_displays7seg_qsys_inst_displays7seg_external_interface_bfm:sig_conduit3
	wire  [6:0] avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit2; // avalon_displays7seg_qsys_inst:displays7seg_external_interface_conduit2 -> avalon_displays7seg_qsys_inst_displays7seg_external_interface_bfm:sig_conduit2
	wire  [6:0] avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit5; // avalon_displays7seg_qsys_inst:displays7seg_external_interface_conduit5 -> avalon_displays7seg_qsys_inst_displays7seg_external_interface_bfm:sig_conduit5
	wire  [6:0] avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit4; // avalon_displays7seg_qsys_inst:displays7seg_external_interface_conduit4 -> avalon_displays7seg_qsys_inst_displays7seg_external_interface_bfm:sig_conduit4
	wire  [6:0] avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit1; // avalon_displays7seg_qsys_inst:displays7seg_external_interface_conduit1 -> avalon_displays7seg_qsys_inst_displays7seg_external_interface_bfm:sig_conduit1
	wire  [6:0] avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit0; // avalon_displays7seg_qsys_inst:displays7seg_external_interface_conduit0 -> avalon_displays7seg_qsys_inst_displays7seg_external_interface_bfm:sig_conduit0
	wire  [6:0] avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit7; // avalon_displays7seg_qsys_inst:displays7seg_external_interface_conduit7 -> avalon_displays7seg_qsys_inst_displays7seg_external_interface_bfm:sig_conduit7
	wire  [6:0] avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit6; // avalon_displays7seg_qsys_inst:displays7seg_external_interface_conduit6 -> avalon_displays7seg_qsys_inst_displays7seg_external_interface_bfm:sig_conduit6
	wire        avalon_displays7seg_qsys_inst_reset_bfm_reset_reset;                    // avalon_displays7seg_qsys_inst_reset_bfm:reset -> [avalon_displays7seg_qsys_inst:reset_reset_n, avalon_displays7seg_qsys_inst_displays7seg_external_interface_bfm:reset]

	avalon_displays7seg_qsys avalon_displays7seg_qsys_inst (
		.clk_clk                                  (avalon_displays7seg_qsys_inst_clk_bfm_clk_clk),                          //                             clk.clk
		.displays7seg_external_interface_conduit0 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit0), // displays7seg_external_interface.conduit0
		.displays7seg_external_interface_conduit1 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit1), //                                .conduit1
		.displays7seg_external_interface_conduit2 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit2), //                                .conduit2
		.displays7seg_external_interface_conduit3 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit3), //                                .conduit3
		.displays7seg_external_interface_conduit4 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit4), //                                .conduit4
		.displays7seg_external_interface_conduit5 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit5), //                                .conduit5
		.displays7seg_external_interface_conduit6 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit6), //                                .conduit6
		.displays7seg_external_interface_conduit7 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit7), //                                .conduit7
		.reset_reset_n                            (avalon_displays7seg_qsys_inst_reset_bfm_reset_reset)                     //                           reset.reset_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) avalon_displays7seg_qsys_inst_clk_bfm (
		.clk (avalon_displays7seg_qsys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm avalon_displays7seg_qsys_inst_displays7seg_external_interface_bfm (
		.clk          (avalon_displays7seg_qsys_inst_clk_bfm_clk_clk),                          //     clk.clk
		.reset        (~avalon_displays7seg_qsys_inst_reset_bfm_reset_reset),                   //   reset.reset
		.sig_conduit0 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit0), // conduit.conduit0
		.sig_conduit1 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit1), //        .conduit1
		.sig_conduit2 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit2), //        .conduit2
		.sig_conduit3 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit3), //        .conduit3
		.sig_conduit4 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit4), //        .conduit4
		.sig_conduit5 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit5), //        .conduit5
		.sig_conduit6 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit6), //        .conduit6
		.sig_conduit7 (avalon_displays7seg_qsys_inst_displays7seg_external_interface_conduit7)  //        .conduit7
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) avalon_displays7seg_qsys_inst_reset_bfm (
		.reset (avalon_displays7seg_qsys_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (avalon_displays7seg_qsys_inst_clk_bfm_clk_clk)        //   clk.clk
	);

endmodule
